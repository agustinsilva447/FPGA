library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ej7a is
port( clk, din: in std_logic;
				 f: out std_logic
);
end ej7a;

architecture hdlc of ej7a is
begin
	
end hdlc;